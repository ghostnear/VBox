module emulator_gameboy

pub struct Config {
	rom_path  string
	bios_path string
}
