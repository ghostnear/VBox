module locale

const map_ro = {
	"language_name": "Română"
	"info_log_app_version": "Versiune: "
	"info_log_session_info": "Informație despre sesiune:"
	"info_log_compiled_with": "Compilat folosind "
	"info_log_language_name": "Limba: "
	"info_log_exit_properly": "Aplicația s-a încheiat cu success."
	"info_log_init_properly": "Aplicația a fost inițializată cu success."
	"message_check_logfile": "Verifică log-ul din folderul executabilului pentru mai multe informații."
	"message_fatal_error_title": "Eroare fatală: "
	"message_unknown_graphics_selected": "Mod de display necunoscut!"
	"message_sdl_could_not_create_window": "Nu a putut fi creată fereastra folosind SDL!"
	"message_sdl_could_not_create_renderer": "Nu a putut fi creat renderer-ul folosind SDL!"
}