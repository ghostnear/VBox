module emulator_gameboy

pub struct Config {
}
