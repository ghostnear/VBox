module chip8

[heap]
struct Timers
{

}