module chip8

// TODO: replace this with a binary file and using the $embed_file() preprocessor.

const font_lowres = [
	u8(0xF0),
	0x90,
	0x90,
	0x90,
	0xF0
	// 0
	0x20,
	0x60,
	0x20,
	0x20,
	0x70
	// 1
	0xF0,
	0x10,
	0xF0,
	0x80,
	0xF0
	// 2
	0xF0,
	0x10,
	0xF0,
	0x10,
	0xF0
	// 3
	0x90,
	0x90,
	0xF0,
	0x10,
	0x10
	// 4
	0xF0,
	0x80,
	0xF0,
	0x10,
	0xF0
	// 5
	0xF0,
	0x80,
	0xF0,
	0x90,
	0xF0
	// 6
	0xF0,
	0x10,
	0x20,
	0x40,
	0x40
	// 7
	0xF0,
	0x90,
	0xF0,
	0x90,
	0xF0
	// 8
	0xF0,
	0x90,
	0xF0,
	0x10,
	0xF0
	// 9
	0xF0,
	0x90,
	0xF0,
	0x90,
	0x90
	// A
	0xE0,
	0x90,
	0xE0,
	0x90,
	0xE0
	// B
	0xF0,
	0x80,
	0x80,
	0x80,
	0xF0
	// C
	0xE0,
	0x90,
	0x90,
	0x90,
	0xE0
	// D
	0xF0,
	0x80,
	0xF0,
	0x80,
	0xF0
	// E
	0xF0,
	0x80,
	0xF0,
	0x80,
	0x80
	// F
]

const font_highres = [
	u8(0xff),
	0xff,
	0xc3,
	0xc3,
	0xc3,
	0xc3,
	0xc3,
	0xc3,
	0xff,
	0xff
	// 0
	0x0c,
	0x0c,
	0x3c,
	0x3c,
	0x0c,
	0x0c,
	0x0c,
	0x0c,
	0x3f,
	0x3f
	// 1
	0xff,
	0xff,
	0x03,
	0x03,
	0xff,
	0xff,
	0xc0,
	0xc0,
	0xff,
	0xff
	// 2
	0xff,
	0xff,
	0x03,
	0x03,
	0xff,
	0xff,
	0x03,
	0x03,
	0xff,
	0xff
	// 3
	0xc3,
	0xc3,
	0xc3,
	0xc3,
	0xff,
	0xff,
	0x03,
	0x03,
	0x03,
	0x03
	// 4
	0xff,
	0xff,
	0xc0,
	0xc0,
	0xff,
	0xff,
	0x03,
	0x03,
	0xff,
	0xff
	// 5
	0xff,
	0xff,
	0xc0,
	0xc0,
	0xff,
	0xff,
	0xc3,
	0xc3,
	0xff,
	0xff
	// 6
	0xff,
	0xff,
	0x03,
	0x03,
	0x0c,
	0x0c,
	0x30,
	0x30,
	0x30,
	0x30
	// 7
	0xff,
	0xff,
	0xc3,
	0xc3,
	0xff,
	0xff,
	0xc3,
	0xc3,
	0xff,
	0xff
	// 8
	0xff,
	0xff,
	0xc3,
	0xc3,
	0xff,
	0xff,
	0x03,
	0x03,
	0xff,
	0xff
	// 9
]
