module chip8

[heap]
struct Audio {
	// TODO: soon
}
