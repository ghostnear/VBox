module emulator_chip8

pub struct Config {
	rom_path         string
	instruction_rate f64
}
