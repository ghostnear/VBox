module chip8

struct Input
{

}