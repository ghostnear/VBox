module chip8

struct Timers
{

}