module chip8

struct Display
{

}