module utilities

pub struct Vec2[T] {
pub mut:
	x T
	y T
}
