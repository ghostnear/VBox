module emulator_dummy

pub struct Config {
}
