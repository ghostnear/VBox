module sdl_driver

pub struct WindowConfig {
	width  int
	height int
	title  string
}
