module chip8

[heap]
struct Input
{

}