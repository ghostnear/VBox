module chip8

[heap]
struct Timers
{
pub mut:
	dt u8
	st u8
}