module locale

// Constant map for the English language.
const map_en = {
	'language_name':                         'English'
	'info_log_quitting':                     'Quitting app...'
	'info_log_app_version':                  'App version: %s'
	'info_log_session_info':                 'Information about this session:'
	'info_log_compiled_with':                'Compiled with %s'
	'info_log_language_name':                'Language: %s (%s)'
	'info_log_exit_properly':                'App exited properly.'
	'info_log_init_properly':                'App was initialized properly.'
	'message_check_logfile':                 "Check the log file in the executable's path for more info."
	'message_fatal_error_title':             'Fatal error: %s'
	'message_unknown_graphics_selected':     'Unknown display mode selected!'
	'message_sdl_could_not_create_window':   'Could not create SDL Window!'
	'message_sdl_could_not_create_renderer': 'Could not create SDL Renderer!'
}
