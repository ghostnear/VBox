module core

// TODO: find a way to extract this from the vmod.
pub const app_version_minor = '1'

pub const app_version_middle = '1'

pub const app_version_major = '0'

pub const app_version = '${app_version_major}.${app_version_middle}.${app_version_minor}'
