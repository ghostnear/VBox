module chip8

struct Audio
{

}